library ieee;
use ieee.std_logic_1164.all;

--Entity
Entity Comparator2 is
	generic ( n: integer :=8);--<-- nbits
	Port(
		A: in std_logic_vector(n-1 downto 0);
		B: in std_logic_vector(n-1 downto 0);
		en: in std_logic;
		AmenorB, AmayorB, AigualB: out std_logic);
end Comparator2;

--Architecture
Architecture solve of Comparator2 is
	-- Signals,Constants,Variables,Components
	Begin
		AmenorB<='1' when A<B and en = '1' else '0';
		AmayorB<='1' when A>B and en = '1' else '0';
		AigualB<='1' when A=B and en = '1' else '0';
end solve;